module RegisterFile
   (input  logic [7:0] din,
    input  logic [3:0] addr,
    input  logic clock, reset_L,
    input  logic read, write,   
    output logic [7:0] dout,
    output logic error);

// Put your code here

endmodule : RegisterFile
